* RC step-response test circuit
* Input: 0->5 V pulse
* Nodes: in (step input), out (capacitor voltage), 0 (ground)

VSTEP in 0 PULSE(0 5 0 1u 1u 0.5m 1m)
R1 in out 1k
C1 out 0 1u

.TRAN 10u 5m
.PRINT TRAN V(out)
.END
